module mult(
  input wire [31:0] A,
  input wire [31:0] B,
  output wire [31:0] Hi,
  output wire [31:0] Lo
);

  // booth algorithm

endmodule
